// main program
module (
    
);

endmodule 